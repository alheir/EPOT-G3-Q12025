.subckt sg3525a INV NI SYN OSC CT RT DCH SS CMP SHD OUA GND VC OUB VIN VRF
A1 N017 0 N009 0 0 N017 N020 0 DFLOP Vhigh=5.1 Trise=20n Rout=30
A2 N018 N019 N009 0 N020 N005 N011 0 OR Vhigh=5.1 Trise=400n Rout=30
A3 N017 N009 0 N019 N018 N023 N022 0 OR Vhigh=5.1 Trise=400n Rout=30
S1 OUA N004 N005 0 HOUT
S2 N012 OUA N011 0 LOUT
S3 OUB N021 N023 0 HOUT
S4 N028 OUB N022 0 LOUT
I1 N031 0 21m
D1 0 N031 IDEAL
R1 N029 N031 8.93
R2 N029 0 22.6
D2 N029 N032 D1_75
D3 0 N032 IDEAL
I2 N032 0 188m
R3 N032 0 2.28
D4 N028 N029 IDEAL
I3 N014 0 21m
D5 0 N014 IDEAL
R4 N013 N014 8.93
R5 N013 0 22.6
D6 N013 N015 D1_75
D7 0 N015 IDEAL
I4 N015 0 188m
R6 N015 0 2.28
D8 N012 N013 IDEAL
D9 VC N021 IDEAL
D10 VC N004 IDEAL
G1 0 N024 NI N027 table=(-70m -100u,0 0,70m 100u)
R7 N024 0 4meg
C1 N024 0 100p
R8 N024 CMP 30
R9 INV 0 1meg
R10 NI 0 1meg
I7 0 VRF 80m
R11 VRF 0 170
D11 0 VRF Z5_1
D12 0 VC Z40
A4 VIN 0 0 0 0 N001 0 0 SCHMITT Vhigh=5.1 Vlow=0.45 Trise=20n Vt=7.25 Vh=0.25
I8 VIN 0 TBL(0 0 3 3.8m 7 19m 8 20m 40 24.1m)
D13 N030 N024 Z5_6
V1 N030 0 0.2
R12 N036 0 5k
R13 SHD N002 5k
Q1 SS N002 N036 0 NPN
D14 N002 0 D1_2
R14 N001 N002 60k
D15 0 SS Z5_1
I9 0 SS 50µ
A5 N002 0 0 0 0 0 N019 0 SCHMITT Vhigh=5.1 Trise=400n Vt=634m Vh=1m
A6 N026 N009 0 0 0 0 N018 0 SRFLOP Vhigh=5.1 Trise=20n Rout=30
A7 0 N025 N019 0 0 0 N026 0 OR Vhigh=5.1 Trise=20n Rout=30
A8 CT N034 0 0 0 0 N025 0 SCHMITT Vhigh=5.1 Trise=20n Vt=0 Vh=10m
E1 N033 0 N024 0 1
E2 N035 0 SS 0 1
R15 N033 N034 500
D16 N034 N035 IDEAL
R16 INV N027 1k
C2 NI N027 40p
R17 SYN 0 2k
R18 OSC N016 250
V2 N003 0 3.64
F1 0 CT V2 -1
D17 N003 RT IDEAL
R19 N016 0 3k
D18 N009 N016 D1_6
S5 0 DCH N009 0 LSW
D19 0 CT Z5_1
A9 N008 N010 0 0 0 0 N009 0 SRFLOP Vhigh=5.1 Ref=0.9 Trise=150n Tfall=250n
A10 N006 N007 0 0 0 0 N008 0 OR Vhigh=5.1 Trise=20n
A11 CT 0 0 0 0 0 N006 0 BUF Vhigh=5.1 Ref=3.2 Trise=20n
A12 CT 0 0 0 0 N010 0 0 BUF Vhigh=5.1 Ref=0.9 Trise=20n
A13 SYN 0 0 0 0 0 N007 0 BUF Vhigh=5.1 Ref=2 Trise=20n
.model NPN NPN
.model PNP PNP
.model HOUT SW(Ron=2.7 Roff=175k Vt=2.8 Vh=-2.1 Vser=1.1 Ilimit=0.6)
.model LOUT SW(Ron=10m Roff=175k Vt=2.8 Vh=-2.1 Vser=0 Ilimit=0.6)
.model IDEAL D(Ron=0 Roff=1G Vfwd=0)
.model D1_75 D(Ron=1.57 Roff=1G Vfwd=1.75)
.model D1_6 D(Ron=0 Roff=1G Vfwd=1.6)
.model Z5_1 D(Ron=1 Roff=1G Vrev=5.075)
.model Z40 D(Ron=0 Roff=175k Vrev=40)
.model Z5_6 D(Ron=1 Roff=1G Vrev=5.6)
.model D1_2 D(Ron=0 Roff=1G Vfwd=1.2)
.model LSW SW(Vt=2.55 Vh=-0.5 Ron=50 Roff=1meg Vser=0.3 Ilimit=50ma)
.ends sg3525a
